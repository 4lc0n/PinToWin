** Profile: "SCHEMATIC1-Solenoid_Driver"  [ c:\users\markl\documents\sem7\smartsystems\pintowin\schematics\main_control\main_control_board-pspicefiles\schematic1\solenoid_driver.sim ] 

** Creating circuit file "Solenoid_Driver.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\markl\Documents\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 3m 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
